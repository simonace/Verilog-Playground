//---------------------------------------------------------------------------
// This arbiter can be used to replace the arbiter in the multi-layer
// AHB Bus Matrix offered by ARM System Design Kit. This arbiter appears
// with the same interface/portlist aiming to easy replacement/integration.
// However, an arbitration strategy of combinatorial logic is implemented
// with the advantage of saving one cycle. Namely the arbitration results
// addr_in_port and no_port are available "instantly" within the same
// cycle the requests comes, rather than a cycle delay in the ARM original
// one. The downside is longer combinatorial path to balance, along with a
// bit overheads.
//
// This file is generated by a Python script giving a parameter of the number
// of input ports. The script is authored by Cheng Cai.
//---------------------------------------------------------------------------

`timescale 1ns/1ps

module ArbiterComb_x4(

    input   wire            HCLK        ,
    input   wire            HRESETn     ,

    input   wire            req_port0   ,
    input   wire            req_port1   ,
    input   wire            req_port2   ,
    input   wire            req_port3   ,

    input   wire            HREADYM     ,
    input   wire            HSELM       ,
    input   wire    [1:0]   HTRANSM     ,
    input   wire            HMASTLOCKM  ,

    output  reg     [1:0]   addr_in_port,
    output  wire            no_port     

);

reg     [1:0]   last_addr_in_port;


assign no_port = ~(req_port0 | req_port1 | req_port2 | req_port3) | ~HREADYM;

always @(*) begin
    if (last_addr_in_port==2'd0) begin
        if (req_port1) begin
            addr_in_port = 2'd1;
        end
        else if (req_port2) begin
            addr_in_port = 2'd2;
        end
        else if (req_port3) begin
            addr_in_port = 2'd3;
        end
        else if (req_port0) begin
            addr_in_port = 2'd0;
        end
        else begin
            addr_in_port = 2'd0;
        end
    end
    else if (last_addr_in_port==2'd1) begin
        if (req_port2) begin
            addr_in_port = 2'd2;
        end
        else if (req_port3) begin
            addr_in_port = 2'd3;
        end
        else if (req_port0) begin
            addr_in_port = 2'd0;
        end
        else if (req_port1) begin
            addr_in_port = 2'd1;
        end
        else begin
            addr_in_port = 2'd0;
        end
    end
    else if (last_addr_in_port==2'd2) begin
        if (req_port3) begin
            addr_in_port = 2'd3;
        end
        else if (req_port0) begin
            addr_in_port = 2'd0;
        end
        else if (req_port1) begin
            addr_in_port = 2'd1;
        end
        else if (req_port2) begin
            addr_in_port = 2'd2;
        end
        else begin
            addr_in_port = 2'd0;
        end
    end
    else if (last_addr_in_port==2'd3) begin
        if (req_port0) begin
            addr_in_port = 2'd0;
        end
        else if (req_port1) begin
            addr_in_port = 2'd1;
        end
        else if (req_port2) begin
            addr_in_port = 2'd2;
        end
        else if (req_port3) begin
            addr_in_port = 2'd3;
        end
        else begin
            addr_in_port = 2'd0;
        end
    end
    else begin
        addr_in_port = 2'd0;
    end
end

always @(negedge HRESETn or posedge HCLK) begin
    if (~HRESETn) begin
        last_addr_in_port <= 2'd0;
    end
    else if (~no_port) begin
        last_addr_in_port <= addr_in_port;
    end
end

endmodule
