//---------------------------------------------------------------------------
// This arbiter can be used to replace the arbiter in the multi-layer
// AHB Bus Matrix offered by ARM System Design Kit. This arbiter appears
// with the same interface/portlist aiming to easy replacement/integration.
// However, an arbitration strategy of combinatorial logic is implemented
// with the advantage of saving one cycle. Namely the arbitration results
// addr_in_port and no_port are available "instantly" within the same
// cycle the requests comes, rather than a cycle delay in the ARM original
// one. The downside is longer combinatorial path to balance, along with a
// bit overheads.
//
// This file is generated by a Python script giving a parameter of the number
// of input ports. The script is authored by Cheng Cai.
//---------------------------------------------------------------------------

`timescale 1ns/1ps

module ArbiterComb_x4(

    input   wire            HCLK        ,
    input   wire            HRESETn     ,

    input   wire            req_port0   ,
    input   wire            req_port1   ,
    input   wire            req_port2   ,
    input   wire            req_port3   ,

    input   wire            HREADYM     ,
    input   wire            HSELM       ,
    input   wire    [1:0]   HTRANSM     ,
    input   wire            HMASTLOCKM  ,

    output  reg     [1:0]   addr_in_port,
    output  wire            no_port     

);

wire    no_pend     ;
reg     pend_port0  ;
reg     pend_port1  ;
reg     pend_port2  ;
reg     pend_port3  ;
reg     req_grant0  ;
reg     req_grant1  ;
reg     req_grant2  ;
reg     req_grant3  ;


assign no_port = ~(req_port0 | req_port1 | req_port2 | req_port3 | pend_port0 | pend_port1 | pend_port2 | pend_port3);
assign no_pend = ~(pend_port0 | pend_port1 | pend_port2 | pend_port3);

always @(*) begin
    if (HSELM & (HTRANSM != 2'b00)) begin
        if (pend_port0) begin
            addr_in_port = 2'd0;
            req_grant0 = 1'b0;
            req_grant1 = 1'b0;
            req_grant2 = 1'b0;
            req_grant3 = 1'b0;
        end
        else if (pend_port1) begin
            addr_in_port = 2'd1;
            req_grant0 = 1'b0;
            req_grant1 = 1'b0;
            req_grant2 = 1'b0;
            req_grant3 = 1'b0;
        end
        else if (pend_port2) begin
            addr_in_port = 2'd2;
            req_grant0 = 1'b0;
            req_grant1 = 1'b0;
            req_grant2 = 1'b0;
            req_grant3 = 1'b0;
        end
        else if (pend_port3) begin
            addr_in_port = 2'd3;
            req_grant0 = 1'b0;
            req_grant1 = 1'b0;
            req_grant2 = 1'b0;
            req_grant3 = 1'b0;
        end
        else if (req_port0) begin
            addr_in_port = 2'd0;
            req_grant0 = 1'b1;
            req_grant1 = 1'b0;
            req_grant2 = 1'b0;
            req_grant3 = 1'b0;
        end
        else if (req_port1) begin
            addr_in_port = 2'd1;
            req_grant0 = 1'b0;
            req_grant1 = 1'b1;
            req_grant2 = 1'b0;
            req_grant3 = 1'b0;
        end
        else if (req_port2) begin
            addr_in_port = 2'd2;
            req_grant0 = 1'b0;
            req_grant1 = 1'b0;
            req_grant2 = 1'b1;
            req_grant3 = 1'b0;
        end
        else if (req_port3) begin
            addr_in_port = 2'd3;
            req_grant0 = 1'b0;
            req_grant1 = 1'b0;
            req_grant2 = 1'b0;
            req_grant3 = 1'b1;
        end
        else begin
            addr_in_port = 2'd0;
            req_grant0 = 1'b0;
            req_grant1 = 1'b0;
            req_grant2 = 1'b0;
            req_grant3 = 1'b0;
        end
        end
    end
    else begin
        addr_in_port = 2'd0;
        req_grant0 = 1'b0;
        req_grant1 = 1'b0;
        req_grant2 = 1'b0;
        req_grant3 = 1'b0;
        end
    end
end

always @(negedge HRESETn or posedge HCLK) begin
    if (~HRESETn) begin
        pend_port0 <= 1'b0;
        pend_port1 <= 1'b0;
        pend_port2 <= 1'b0;
        pend_port3 <= 1'b0;
    end
    else begin
        if (~HMASTLOCK & HREADYM) begin
            if (no_pend) begin
                pend_port0 <= ~req_grant0 & req_port0;
                pend_port1 <= ~req_grant1 & req_port1;
                pend_port2 <= ~req_grant2 & req_port2;
                pend_port3 <= ~req_grant3 & req_port3;
            end
            else if (pend_port0) begin
                pend_port0 <= 1'b0;
                pend_port1 <= pend_port1;
                pend_port2 <= pend_port2;
                pend_port3 <= pend_port3;
            end
            else if (pend_port1) begin
                pend_port0 <= 1'b0;
                pend_port1 <= 1'b0;
                pend_port2 <= pend_port2;
                pend_port3 <= pend_port3;
            end
            else if (pend_port2) begin
                pend_port0 <= 1'b0;
                pend_port1 <= 1'b0;
                pend_port2 <= 1'b0;
                pend_port3 <= pend_port3;
            end
            else if (pend_port3) begin
                pend_port0 <= 1'b0;
                pend_port1 <= 1'b0;
                pend_port2 <= 1'b0;
                pend_port3 <= 1'b0;
            end
        end
    end
end

endmodule